// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_proj_example
 *
 * This is an example of a (trivially simple) user project,
 * showing how the user project can connect to the logic
 * analyzer, the wishbone bus, and the I/O pads.
 *
 * This project generates an integer count, which is output
 * on the user area GPIO pads (digital output only).  The
 * wishbone connection allows the project to be controlled
 * (start and stop) from the management SoC program.
 *
 * See the testbenches in directory "mprj_counter" for the
 * example programs that drive this user project.  The three
 * testbenches are "io_ports", "la_test1", and "la_test2".
 *
 *-------------------------------------------------------------
 */

module user_proj_example #(
    parameter BITS = 16
)(
`ifdef USE_POWER_PINS
    inout vdd,	// User area 1 1.8V supply
    inout vss,	// User area 1 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o
);
    wire [31:0] dat_w;
    wire [31:0] dat_r;
    wire sel;
    wire we;
    wire cyc;
    wire stb;
    wire ack;
    wire clk;
    wire rst;
    wire [31:0] adr;
    
    assign dat_w = wbs_dat_i;
    assign wbs_dat_o = dat_r;
    assign sel = wbs_sel_i[0];
    assign we = wbs_we_i;
    assign cyc = wbs_cyc_i;
    assign stb = wbs_stb_i;
    assign wbs_ack_o = ack;
    assign clk = wb_clk_i;
    assign rst = wb_rst_i;
    assign adr = wbs_adr_i;
    
    systolic_array systolic_array(
        .dat_w(dat_w),
        .dat_r(dat_r),
        .sel(sel),
        .we(we),
        .cyc(cyc),
        .stb(stb),
        .ack(ack),
        .clk(clk),
        .rst(rst),
        .adr(adr)
    );

endmodule
 
module systolic_array(dat_w, dat_r, sel, we, cyc, stb, ack, clk, rst, adr);
  reg \$auto$verilog_backend.cc:2097:dump_module$1  = 0;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$103 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$108 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$113 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$118 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$123 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$128 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$13 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$133 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$138 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$143 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$148 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$153 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$158 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$163 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$168 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$173 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$178 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$18 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$183 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$188 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$193 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$198 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$203 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$208 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$213 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$218 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$223 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$228 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$23 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$233 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$238 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$243 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$248 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$253 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$258 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$263 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$268 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$273 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$278 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$28 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$283 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$288 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$293 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$298 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$3 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$303 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$308 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$313 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$318 ;
  (* src = "/home/james/systolicArray.py:34" *)
  wire \$320 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$33 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$38 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$43 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$48 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$53 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$58 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$63 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$68 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$73 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$78 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$8 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$83 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$88 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$93 ;
  (* src = "/home/james/systolicArray.py:21" *)
  wire [31:0] \$98 ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal  = 32'd0;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$1  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$1$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$10  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$10$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$100  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$100$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$101  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$101$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$102  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$102$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$105  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$105$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$106  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$106$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$107  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$107$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$11  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$11$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$110  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$110$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$111  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$111$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$112  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$112$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$115  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$115$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$116  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$116$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$117  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$117$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$12  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$12$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$120  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$120$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$121  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$121$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$122  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$122$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$125  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$125$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$126  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$126$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$127  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$127$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$130  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$130$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$131  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$131$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$132  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$132$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$135  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$135$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$136  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$136$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$137  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$137$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$140  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$140$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$141  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$141$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$142  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$142$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$145  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$145$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$146  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$146$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$147  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$147$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$15  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$15$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$150  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$150$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$151  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$151$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$152  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$152$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$155  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$155$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$156  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$156$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$157  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$157$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$16  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$16$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$160  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$160$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$161  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$161$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$162  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$162$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$165  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$165$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$166  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$166$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$167  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$167$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$17  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$17$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$170  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$170$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$171  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$171$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$172  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$172$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$175  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$175$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$176  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$176$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$177  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$177$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$180  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$180$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$181  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$181$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$182  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$182$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$185  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$185$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$186  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$186$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$187  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$187$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$190  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$190$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$191  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$191$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$192  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$192$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$195  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$195$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$196  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$196$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$197  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$197$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$2  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$2$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$20  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$20$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$200  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$200$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$201  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$201$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$202  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$202$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$205  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$205$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$206  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$206$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$207  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$207$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$21  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$21$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$210  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$210$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$211  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$211$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$212  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$212$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$215  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$215$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$216  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$216$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$217  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$217$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$22  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$22$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$220  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$220$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$221  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$221$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$222  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$222$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$225  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$225$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$226  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$226$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$227  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$227$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$230  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$230$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$231  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$231$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$232  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$232$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$235  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$235$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$236  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$236$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$237  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$237$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$240  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$240$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$241  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$241$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$242  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$242$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$245  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$245$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$246  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$246$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$247  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$247$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$25  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$25$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$250  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$250$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$251  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$251$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$252  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$252$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$255  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$255$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$256  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$256$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$257  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$257$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$26  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$26$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$260  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$260$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$261  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$261$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$262  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$262$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$265  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$265$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$266  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$266$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$267  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$267$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$27  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$27$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$270  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$270$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$271  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$271$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$272  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$272$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$275  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$275$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$276  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$276$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$277  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$277$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$280  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$280$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$281  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$281$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$282  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$282$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$285  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$285$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$286  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$286$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$287  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$287$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$290  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$290$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$291  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$291$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$292  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$292$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$295  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$295$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$296  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$296$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$297  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$297$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$30  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$30$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$300  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$300$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$301  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$301$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$302  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$302$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$305  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$305$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$306  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$306$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$307  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$307$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$31  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$31$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$310  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$310$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$311  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$311$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$312  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$312$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$315  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$315$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$316  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$316$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$317  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$317$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$32  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$32$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$35  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$35$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$36  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$36$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$37  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$37$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$40  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$40$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$41  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$41$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$42  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$42$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$45  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$45$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$46  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$46$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$47  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$47$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$5  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$5$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$50  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$50$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$51  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$51$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$52  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$52$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$55  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$55$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$56  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$56$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$57  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$57$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$6  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$6$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$60  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$60$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$61  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$61$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$62  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$62$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$65  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$65$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$66  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$66$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$67  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$67$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$7  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$7$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$70  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$70$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$71  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$71$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$72  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$72$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$75  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$75$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$76  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$76$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$77  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$77$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$80  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$80$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$81  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$81$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$82  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$82$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$85  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$85$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$86  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$86$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$87  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$87$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$90  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$90$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$91  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$91$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$92  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$92$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$95  = 32'd0;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$95$next ;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$96  = 16'h0000;
  (* src = "/home/james/systolicArray.py:11" *)
  reg [15:0] \$signal$96$next ;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$97  = 16'h0000;
  (* src = "/home/james/systolicArray.py:12" *)
  reg [15:0] \$signal$97$next ;
  (* src = "/home/james/systolicArray.py:13" *)
  reg [31:0] \$signal$next ;
  (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/lib/wiring.py:227" *)
  output ack;
  reg ack = 1'h0;
  (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/lib/wiring.py:227" *)
  reg \ack$next ;
  (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/lib/wiring.py:227" *)
  input [31:0] adr;
  wire [31:0] adr;
  (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/ir.py:508" *)
  input clk;
  wire clk;
  (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/lib/wiring.py:227" *)
  input cyc;
  wire cyc;
  (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/lib/wiring.py:227" *)
  output [31:0] dat_r;
  reg [31:0] dat_r;
  (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/lib/wiring.py:227" *)
  input [31:0] dat_w;
  wire [31:0] dat_w;
  (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/ir.py:508" *)
  input rst;
  wire rst;
  (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/lib/wiring.py:227" *)
  input sel;
  wire sel;
  (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/lib/wiring.py:227" *)
  input stb;
  wire stb;
  (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/lib/wiring.py:227" *)
  input we;
  wire we;
  assign \$103  = \$signal$101  * (* src = "/home/james/systolicArray.py:21" *) \$signal$102 ;
  assign \$108  = \$signal$106  * (* src = "/home/james/systolicArray.py:21" *) \$signal$107 ;
  assign \$113  = \$signal$111  * (* src = "/home/james/systolicArray.py:21" *) \$signal$112 ;
  assign \$118  = \$signal$116  * (* src = "/home/james/systolicArray.py:21" *) \$signal$117 ;
  assign \$123  = \$signal$121  * (* src = "/home/james/systolicArray.py:21" *) \$signal$122 ;
  assign \$128  = \$signal$126  * (* src = "/home/james/systolicArray.py:21" *) \$signal$127 ;
  assign \$133  = \$signal$131  * (* src = "/home/james/systolicArray.py:21" *) \$signal$132 ;
  assign \$138  = \$signal$136  * (* src = "/home/james/systolicArray.py:21" *) \$signal$137 ;
  assign \$13  = \$signal$11  * (* src = "/home/james/systolicArray.py:21" *) \$signal$12 ;
  assign \$143  = \$signal$141  * (* src = "/home/james/systolicArray.py:21" *) \$signal$142 ;
  assign \$148  = \$signal$146  * (* src = "/home/james/systolicArray.py:21" *) \$signal$147 ;
  assign \$153  = \$signal$151  * (* src = "/home/james/systolicArray.py:21" *) \$signal$152 ;
  assign \$158  = \$signal$156  * (* src = "/home/james/systolicArray.py:21" *) \$signal$157 ;
  assign \$163  = \$signal$161  * (* src = "/home/james/systolicArray.py:21" *) \$signal$162 ;
  assign \$168  = \$signal$166  * (* src = "/home/james/systolicArray.py:21" *) \$signal$167 ;
  assign \$173  = \$signal$171  * (* src = "/home/james/systolicArray.py:21" *) \$signal$172 ;
  assign \$178  = \$signal$176  * (* src = "/home/james/systolicArray.py:21" *) \$signal$177 ;
  assign \$183  = \$signal$181  * (* src = "/home/james/systolicArray.py:21" *) \$signal$182 ;
  assign \$188  = \$signal$186  * (* src = "/home/james/systolicArray.py:21" *) \$signal$187 ;
  assign \$18  = \$signal$16  * (* src = "/home/james/systolicArray.py:21" *) \$signal$17 ;
  assign \$193  = \$signal$191  * (* src = "/home/james/systolicArray.py:21" *) \$signal$192 ;
  assign \$198  = \$signal$196  * (* src = "/home/james/systolicArray.py:21" *) \$signal$197 ;
  assign \$203  = \$signal$201  * (* src = "/home/james/systolicArray.py:21" *) \$signal$202 ;
  assign \$208  = \$signal$206  * (* src = "/home/james/systolicArray.py:21" *) \$signal$207 ;
  assign \$213  = \$signal$211  * (* src = "/home/james/systolicArray.py:21" *) \$signal$212 ;
  assign \$218  = \$signal$216  * (* src = "/home/james/systolicArray.py:21" *) \$signal$217 ;
  assign \$223  = \$signal$221  * (* src = "/home/james/systolicArray.py:21" *) \$signal$222 ;
  assign \$228  = \$signal$226  * (* src = "/home/james/systolicArray.py:21" *) \$signal$227 ;
  assign \$233  = \$signal$231  * (* src = "/home/james/systolicArray.py:21" *) \$signal$232 ;
  assign \$238  = \$signal$236  * (* src = "/home/james/systolicArray.py:21" *) \$signal$237 ;
  assign \$23  = \$signal$21  * (* src = "/home/james/systolicArray.py:21" *) \$signal$22 ;
  assign \$243  = \$signal$241  * (* src = "/home/james/systolicArray.py:21" *) \$signal$242 ;
  assign \$248  = \$signal$246  * (* src = "/home/james/systolicArray.py:21" *) \$signal$247 ;
  assign \$253  = \$signal$251  * (* src = "/home/james/systolicArray.py:21" *) \$signal$252 ;
  assign \$258  = \$signal$256  * (* src = "/home/james/systolicArray.py:21" *) \$signal$257 ;
  assign \$263  = \$signal$261  * (* src = "/home/james/systolicArray.py:21" *) \$signal$262 ;
  assign \$268  = \$signal$266  * (* src = "/home/james/systolicArray.py:21" *) \$signal$267 ;
  assign \$273  = \$signal$271  * (* src = "/home/james/systolicArray.py:21" *) \$signal$272 ;
  assign \$278  = \$signal$276  * (* src = "/home/james/systolicArray.py:21" *) \$signal$277 ;
  assign \$283  = \$signal$281  * (* src = "/home/james/systolicArray.py:21" *) \$signal$282 ;
  assign \$288  = \$signal$286  * (* src = "/home/james/systolicArray.py:21" *) \$signal$287 ;
  assign \$28  = \$signal$26  * (* src = "/home/james/systolicArray.py:21" *) \$signal$27 ;
  assign \$293  = \$signal$291  * (* src = "/home/james/systolicArray.py:21" *) \$signal$292 ;
  assign \$298  = \$signal$296  * (* src = "/home/james/systolicArray.py:21" *) \$signal$297 ;
  assign \$303  = \$signal$301  * (* src = "/home/james/systolicArray.py:21" *) \$signal$302 ;
  assign \$308  = \$signal$306  * (* src = "/home/james/systolicArray.py:21" *) \$signal$307 ;
  assign \$313  = \$signal$311  * (* src = "/home/james/systolicArray.py:21" *) \$signal$312 ;
  assign \$318  = \$signal$316  * (* src = "/home/james/systolicArray.py:21" *) \$signal$317 ;
  assign \$320  = cyc & (* src = "/home/james/systolicArray.py:34" *) stb;
  always @(posedge clk)
    \$signal  <= \$signal$next ;
  always @(posedge clk)
    \$signal$5  <= \$signal$5$next ;
  always @(posedge clk)
    \$signal$10  <= \$signal$10$next ;
  always @(posedge clk)
    \$signal$15  <= \$signal$15$next ;
  always @(posedge clk)
    \$signal$20  <= \$signal$20$next ;
  always @(posedge clk)
    \$signal$25  <= \$signal$25$next ;
  always @(posedge clk)
    \$signal$30  <= \$signal$30$next ;
  always @(posedge clk)
    \$signal$35  <= \$signal$35$next ;
  always @(posedge clk)
    \$signal$40  <= \$signal$40$next ;
  always @(posedge clk)
    \$signal$45  <= \$signal$45$next ;
  always @(posedge clk)
    \$signal$50  <= \$signal$50$next ;
  always @(posedge clk)
    \$signal$55  <= \$signal$55$next ;
  always @(posedge clk)
    \$signal$60  <= \$signal$60$next ;
  always @(posedge clk)
    \$signal$65  <= \$signal$65$next ;
  always @(posedge clk)
    \$signal$70  <= \$signal$70$next ;
  always @(posedge clk)
    \$signal$75  <= \$signal$75$next ;
  always @(posedge clk)
    \$signal$80  <= \$signal$80$next ;
  always @(posedge clk)
    \$signal$85  <= \$signal$85$next ;
  assign \$33  = \$signal$31  * (* src = "/home/james/systolicArray.py:21" *) \$signal$32 ;
  always @(posedge clk)
    \$signal$90  <= \$signal$90$next ;
  always @(posedge clk)
    \$signal$95  <= \$signal$95$next ;
  always @(posedge clk)
    \$signal$100  <= \$signal$100$next ;
  always @(posedge clk)
    \$signal$105  <= \$signal$105$next ;
  always @(posedge clk)
    \$signal$110  <= \$signal$110$next ;
  always @(posedge clk)
    \$signal$115  <= \$signal$115$next ;
  always @(posedge clk)
    \$signal$120  <= \$signal$120$next ;
  always @(posedge clk)
    \$signal$125  <= \$signal$125$next ;
  always @(posedge clk)
    \$signal$130  <= \$signal$130$next ;
  always @(posedge clk)
    \$signal$135  <= \$signal$135$next ;
  always @(posedge clk)
    \$signal$140  <= \$signal$140$next ;
  always @(posedge clk)
    \$signal$145  <= \$signal$145$next ;
  always @(posedge clk)
    \$signal$150  <= \$signal$150$next ;
  always @(posedge clk)
    \$signal$155  <= \$signal$155$next ;
  always @(posedge clk)
    \$signal$160  <= \$signal$160$next ;
  always @(posedge clk)
    \$signal$165  <= \$signal$165$next ;
  always @(posedge clk)
    \$signal$170  <= \$signal$170$next ;
  always @(posedge clk)
    \$signal$175  <= \$signal$175$next ;
  always @(posedge clk)
    \$signal$180  <= \$signal$180$next ;
  always @(posedge clk)
    \$signal$185  <= \$signal$185$next ;
  always @(posedge clk)
    \$signal$190  <= \$signal$190$next ;
  always @(posedge clk)
    \$signal$195  <= \$signal$195$next ;
  always @(posedge clk)
    \$signal$200  <= \$signal$200$next ;
  always @(posedge clk)
    \$signal$205  <= \$signal$205$next ;
  always @(posedge clk)
    \$signal$210  <= \$signal$210$next ;
  always @(posedge clk)
    \$signal$215  <= \$signal$215$next ;
  always @(posedge clk)
    \$signal$220  <= \$signal$220$next ;
  always @(posedge clk)
    \$signal$225  <= \$signal$225$next ;
  always @(posedge clk)
    \$signal$230  <= \$signal$230$next ;
  always @(posedge clk)
    \$signal$235  <= \$signal$235$next ;
  always @(posedge clk)
    \$signal$240  <= \$signal$240$next ;
  always @(posedge clk)
    \$signal$245  <= \$signal$245$next ;
  always @(posedge clk)
    \$signal$250  <= \$signal$250$next ;
  always @(posedge clk)
    \$signal$255  <= \$signal$255$next ;
  always @(posedge clk)
    \$signal$260  <= \$signal$260$next ;
  always @(posedge clk)
    \$signal$265  <= \$signal$265$next ;
  always @(posedge clk)
    \$signal$270  <= \$signal$270$next ;
  always @(posedge clk)
    \$signal$275  <= \$signal$275$next ;
  always @(posedge clk)
    \$signal$280  <= \$signal$280$next ;
  always @(posedge clk)
    \$signal$285  <= \$signal$285$next ;
  always @(posedge clk)
    \$signal$290  <= \$signal$290$next ;
  always @(posedge clk)
    \$signal$295  <= \$signal$295$next ;
  always @(posedge clk)
    \$signal$300  <= \$signal$300$next ;
  always @(posedge clk)
    \$signal$305  <= \$signal$305$next ;
  always @(posedge clk)
    \$signal$310  <= \$signal$310$next ;
  always @(posedge clk)
    \$signal$315  <= \$signal$315$next ;
  always @(posedge clk)
    \$signal$1  <= \$signal$1$next ;
  always @(posedge clk)
    \$signal$2  <= \$signal$2$next ;
  always @(posedge clk)
    \$signal$6  <= \$signal$6$next ;
  always @(posedge clk)
    \$signal$7  <= \$signal$7$next ;
  assign \$38  = \$signal$36  * (* src = "/home/james/systolicArray.py:21" *) \$signal$37 ;
  always @(posedge clk)
    \$signal$11  <= \$signal$11$next ;
  always @(posedge clk)
    \$signal$12  <= \$signal$12$next ;
  always @(posedge clk)
    \$signal$16  <= \$signal$16$next ;
  always @(posedge clk)
    \$signal$17  <= \$signal$17$next ;
  always @(posedge clk)
    \$signal$21  <= \$signal$21$next ;
  always @(posedge clk)
    \$signal$22  <= \$signal$22$next ;
  always @(posedge clk)
    \$signal$26  <= \$signal$26$next ;
  always @(posedge clk)
    \$signal$27  <= \$signal$27$next ;
  always @(posedge clk)
    \$signal$31  <= \$signal$31$next ;
  always @(posedge clk)
    \$signal$32  <= \$signal$32$next ;
  assign \$3  = \$signal$1  * (* src = "/home/james/systolicArray.py:21" *) \$signal$2 ;
  always @(posedge clk)
    \$signal$36  <= \$signal$36$next ;
  always @(posedge clk)
    \$signal$37  <= \$signal$37$next ;
  always @(posedge clk)
    \$signal$41  <= \$signal$41$next ;
  always @(posedge clk)
    \$signal$42  <= \$signal$42$next ;
  always @(posedge clk)
    \$signal$46  <= \$signal$46$next ;
  always @(posedge clk)
    \$signal$47  <= \$signal$47$next ;
  always @(posedge clk)
    \$signal$51  <= \$signal$51$next ;
  always @(posedge clk)
    \$signal$52  <= \$signal$52$next ;
  always @(posedge clk)
    \$signal$56  <= \$signal$56$next ;
  always @(posedge clk)
    \$signal$57  <= \$signal$57$next ;
  always @(posedge clk)
    \$signal$61  <= \$signal$61$next ;
  always @(posedge clk)
    \$signal$62  <= \$signal$62$next ;
  always @(posedge clk)
    \$signal$66  <= \$signal$66$next ;
  always @(posedge clk)
    \$signal$67  <= \$signal$67$next ;
  always @(posedge clk)
    \$signal$71  <= \$signal$71$next ;
  always @(posedge clk)
    \$signal$72  <= \$signal$72$next ;
  always @(posedge clk)
    \$signal$76  <= \$signal$76$next ;
  always @(posedge clk)
    \$signal$77  <= \$signal$77$next ;
  always @(posedge clk)
    \$signal$81  <= \$signal$81$next ;
  always @(posedge clk)
    \$signal$82  <= \$signal$82$next ;
  always @(posedge clk)
    \$signal$86  <= \$signal$86$next ;
  always @(posedge clk)
    \$signal$87  <= \$signal$87$next ;
  always @(posedge clk)
    \$signal$91  <= \$signal$91$next ;
  always @(posedge clk)
    \$signal$92  <= \$signal$92$next ;
  always @(posedge clk)
    \$signal$96  <= \$signal$96$next ;
  always @(posedge clk)
    \$signal$97  <= \$signal$97$next ;
  always @(posedge clk)
    \$signal$101  <= \$signal$101$next ;
  always @(posedge clk)
    \$signal$102  <= \$signal$102$next ;
  always @(posedge clk)
    \$signal$106  <= \$signal$106$next ;
  always @(posedge clk)
    \$signal$107  <= \$signal$107$next ;
  always @(posedge clk)
    \$signal$111  <= \$signal$111$next ;
  always @(posedge clk)
    \$signal$112  <= \$signal$112$next ;
  always @(posedge clk)
    \$signal$116  <= \$signal$116$next ;
  always @(posedge clk)
    \$signal$117  <= \$signal$117$next ;
  always @(posedge clk)
    \$signal$121  <= \$signal$121$next ;
  always @(posedge clk)
    \$signal$122  <= \$signal$122$next ;
  always @(posedge clk)
    \$signal$126  <= \$signal$126$next ;
  always @(posedge clk)
    \$signal$127  <= \$signal$127$next ;
  always @(posedge clk)
    \$signal$131  <= \$signal$131$next ;
  always @(posedge clk)
    \$signal$132  <= \$signal$132$next ;
  assign \$43  = \$signal$41  * (* src = "/home/james/systolicArray.py:21" *) \$signal$42 ;
  always @(posedge clk)
    \$signal$136  <= \$signal$136$next ;
  always @(posedge clk)
    \$signal$137  <= \$signal$137$next ;
  always @(posedge clk)
    \$signal$141  <= \$signal$141$next ;
  always @(posedge clk)
    \$signal$142  <= \$signal$142$next ;
  always @(posedge clk)
    \$signal$146  <= \$signal$146$next ;
  always @(posedge clk)
    \$signal$147  <= \$signal$147$next ;
  always @(posedge clk)
    \$signal$151  <= \$signal$151$next ;
  always @(posedge clk)
    \$signal$152  <= \$signal$152$next ;
  always @(posedge clk)
    \$signal$156  <= \$signal$156$next ;
  always @(posedge clk)
    \$signal$157  <= \$signal$157$next ;
  always @(posedge clk)
    \$signal$161  <= \$signal$161$next ;
  always @(posedge clk)
    \$signal$162  <= \$signal$162$next ;
  always @(posedge clk)
    \$signal$166  <= \$signal$166$next ;
  always @(posedge clk)
    \$signal$167  <= \$signal$167$next ;
  always @(posedge clk)
    \$signal$171  <= \$signal$171$next ;
  always @(posedge clk)
    \$signal$172  <= \$signal$172$next ;
  always @(posedge clk)
    \$signal$176  <= \$signal$176$next ;
  always @(posedge clk)
    \$signal$177  <= \$signal$177$next ;
  always @(posedge clk)
    \$signal$181  <= \$signal$181$next ;
  always @(posedge clk)
    \$signal$182  <= \$signal$182$next ;
  always @(posedge clk)
    \$signal$186  <= \$signal$186$next ;
  always @(posedge clk)
    \$signal$187  <= \$signal$187$next ;
  always @(posedge clk)
    \$signal$191  <= \$signal$191$next ;
  always @(posedge clk)
    \$signal$192  <= \$signal$192$next ;
  always @(posedge clk)
    \$signal$196  <= \$signal$196$next ;
  always @(posedge clk)
    \$signal$197  <= \$signal$197$next ;
  always @(posedge clk)
    \$signal$201  <= \$signal$201$next ;
  always @(posedge clk)
    \$signal$202  <= \$signal$202$next ;
  always @(posedge clk)
    \$signal$206  <= \$signal$206$next ;
  always @(posedge clk)
    \$signal$207  <= \$signal$207$next ;
  always @(posedge clk)
    \$signal$211  <= \$signal$211$next ;
  always @(posedge clk)
    \$signal$212  <= \$signal$212$next ;
  always @(posedge clk)
    \$signal$216  <= \$signal$216$next ;
  always @(posedge clk)
    \$signal$217  <= \$signal$217$next ;
  always @(posedge clk)
    \$signal$221  <= \$signal$221$next ;
  always @(posedge clk)
    \$signal$222  <= \$signal$222$next ;
  always @(posedge clk)
    \$signal$226  <= \$signal$226$next ;
  always @(posedge clk)
    \$signal$227  <= \$signal$227$next ;
  always @(posedge clk)
    \$signal$231  <= \$signal$231$next ;
  always @(posedge clk)
    \$signal$232  <= \$signal$232$next ;
  always @(posedge clk)
    \$signal$236  <= \$signal$236$next ;
  always @(posedge clk)
    \$signal$237  <= \$signal$237$next ;
  always @(posedge clk)
    \$signal$241  <= \$signal$241$next ;
  always @(posedge clk)
    \$signal$242  <= \$signal$242$next ;
  always @(posedge clk)
    \$signal$246  <= \$signal$246$next ;
  always @(posedge clk)
    \$signal$247  <= \$signal$247$next ;
  always @(posedge clk)
    \$signal$251  <= \$signal$251$next ;
  always @(posedge clk)
    \$signal$252  <= \$signal$252$next ;
  always @(posedge clk)
    \$signal$256  <= \$signal$256$next ;
  always @(posedge clk)
    \$signal$257  <= \$signal$257$next ;
  assign \$48  = \$signal$46  * (* src = "/home/james/systolicArray.py:21" *) \$signal$47 ;
  always @(posedge clk)
    \$signal$261  <= \$signal$261$next ;
  always @(posedge clk)
    \$signal$262  <= \$signal$262$next ;
  always @(posedge clk)
    \$signal$266  <= \$signal$266$next ;
  always @(posedge clk)
    \$signal$267  <= \$signal$267$next ;
  always @(posedge clk)
    \$signal$271  <= \$signal$271$next ;
  always @(posedge clk)
    \$signal$272  <= \$signal$272$next ;
  always @(posedge clk)
    \$signal$276  <= \$signal$276$next ;
  always @(posedge clk)
    \$signal$277  <= \$signal$277$next ;
  always @(posedge clk)
    \$signal$281  <= \$signal$281$next ;
  always @(posedge clk)
    \$signal$282  <= \$signal$282$next ;
  always @(posedge clk)
    \$signal$286  <= \$signal$286$next ;
  always @(posedge clk)
    \$signal$287  <= \$signal$287$next ;
  always @(posedge clk)
    \$signal$291  <= \$signal$291$next ;
  always @(posedge clk)
    \$signal$292  <= \$signal$292$next ;
  always @(posedge clk)
    \$signal$296  <= \$signal$296$next ;
  always @(posedge clk)
    \$signal$297  <= \$signal$297$next ;
  always @(posedge clk)
    \$signal$301  <= \$signal$301$next ;
  always @(posedge clk)
    \$signal$302  <= \$signal$302$next ;
  always @(posedge clk)
    \$signal$306  <= \$signal$306$next ;
  always @(posedge clk)
    \$signal$307  <= \$signal$307$next ;
  always @(posedge clk)
    \$signal$311  <= \$signal$311$next ;
  always @(posedge clk)
    \$signal$312  <= \$signal$312$next ;
  always @(posedge clk)
    \$signal$316  <= \$signal$316$next ;
  always @(posedge clk)
    \$signal$317  <= \$signal$317$next ;
  always @(posedge clk)
    ack <= \ack$next ;
  assign \$53  = \$signal$51  * (* src = "/home/james/systolicArray.py:21" *) \$signal$52 ;
  assign \$58  = \$signal$56  * (* src = "/home/james/systolicArray.py:21" *) \$signal$57 ;
  assign \$63  = \$signal$61  * (* src = "/home/james/systolicArray.py:21" *) \$signal$62 ;
  assign \$68  = \$signal$66  * (* src = "/home/james/systolicArray.py:21" *) \$signal$67 ;
  assign \$73  = \$signal$71  * (* src = "/home/james/systolicArray.py:21" *) \$signal$72 ;
  assign \$78  = \$signal$76  * (* src = "/home/james/systolicArray.py:21" *) \$signal$77 ;
  assign \$83  = \$signal$81  * (* src = "/home/james/systolicArray.py:21" *) \$signal$82 ;
  assign \$88  = \$signal$86  * (* src = "/home/james/systolicArray.py:21" *) \$signal$87 ;
  assign \$8  = \$signal$6  * (* src = "/home/james/systolicArray.py:21" *) \$signal$7 ;
  assign \$93  = \$signal$91  * (* src = "/home/james/systolicArray.py:21" *) \$signal$92 ;
  assign \$98  = \$signal$96  * (* src = "/home/james/systolicArray.py:21" *) \$signal$97 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$next  = \$3 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$5$next  = \$8 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$5$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$50$next  = \$53 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$50$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$87$next  = \$signal$87 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          \$signal$87$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$87$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$91$next  = \$signal$91 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          \$signal$91$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$91$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$92$next  = \$signal$92 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          \$signal$92$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$92$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$96$next  = \$signal$96 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          \$signal$96$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$96$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$97$next  = \$signal$97 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          \$signal$97$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$97$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$101$next  = \$signal$101 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          \$signal$101$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$101$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$102$next  = \$signal$102 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          \$signal$102$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$102$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$106$next  = \$signal$106 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          \$signal$106$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$106$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$107$next  = \$signal$107 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          \$signal$107$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$107$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$111$next  = \$signal$111 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          \$signal$111$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$111$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$55$next  = \$58 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$55$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$112$next  = \$signal$112 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          \$signal$112$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$112$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$116$next  = \$signal$116 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          \$signal$116$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$116$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$117$next  = \$signal$117 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          \$signal$117$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$117$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$121$next  = \$signal$121 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          \$signal$121$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$121$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$122$next  = \$signal$122 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          \$signal$122$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$122$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$126$next  = \$signal$126 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          \$signal$126$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$126$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$127$next  = \$signal$127 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          \$signal$127$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$127$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$131$next  = \$signal$131 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          \$signal$131$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$131$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$132$next  = \$signal$132 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          \$signal$132$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$132$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$136$next  = \$signal$136 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          \$signal$136$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$136$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$60$next  = \$63 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$60$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$137$next  = \$signal$137 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          \$signal$137$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$137$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$141$next  = \$signal$141 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          \$signal$141$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$141$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$142$next  = \$signal$142 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          \$signal$142$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$142$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$146$next  = \$signal$146 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          \$signal$146$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$146$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$147$next  = \$signal$147 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          \$signal$147$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$147$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$151$next  = \$signal$151 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          \$signal$151$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$151$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$152$next  = \$signal$152 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          \$signal$152$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$152$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$156$next  = \$signal$156 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          \$signal$156$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$156$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$157$next  = \$signal$157 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          \$signal$157$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$157$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$161$next  = \$signal$161 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          \$signal$161$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$161$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$65$next  = \$68 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$65$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$162$next  = \$signal$162 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          \$signal$162$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$162$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$166$next  = \$signal$166 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          \$signal$166$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$166$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$167$next  = \$signal$167 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          \$signal$167$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$167$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$171$next  = \$signal$171 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          \$signal$171$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$171$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$172$next  = \$signal$172 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          \$signal$172$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$172$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$176$next  = \$signal$176 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          \$signal$176$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$176$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$177$next  = \$signal$177 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          \$signal$177$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$177$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$181$next  = \$signal$181 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          \$signal$181$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$181$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$182$next  = \$signal$182 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          \$signal$182$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$182$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$186$next  = \$signal$186 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          \$signal$186$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$186$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$70$next  = \$73 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$70$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$187$next  = \$signal$187 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          \$signal$187$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$187$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$191$next  = \$signal$191 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          \$signal$191$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$191$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$192$next  = \$signal$192 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          \$signal$192$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$192$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$196$next  = \$signal$196 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          \$signal$196$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$196$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$197$next  = \$signal$197 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          \$signal$197$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$197$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$201$next  = \$signal$201 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          \$signal$201$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$201$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$202$next  = \$signal$202 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          \$signal$202$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$202$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$206$next  = \$signal$206 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          \$signal$206$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$206$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$207$next  = \$signal$207 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          \$signal$207$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$207$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$211$next  = \$signal$211 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          \$signal$211$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$211$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$75$next  = \$78 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$75$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$212$next  = \$signal$212 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          \$signal$212$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$212$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$216$next  = \$signal$216 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          \$signal$216$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$216$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$217$next  = \$signal$217 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          \$signal$217$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$217$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$221$next  = \$signal$221 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          \$signal$221$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$221$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$222$next  = \$signal$222 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          \$signal$222$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$222$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$226$next  = \$signal$226 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          \$signal$226$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$226$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$227$next  = \$signal$227 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          \$signal$227$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$227$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$231$next  = \$signal$231 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          \$signal$231$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$231$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$232$next  = \$signal$232 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          \$signal$232$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$232$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$236$next  = \$signal$236 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          \$signal$236$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$236$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$80$next  = \$83 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$80$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$237$next  = \$signal$237 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          \$signal$237$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$237$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$241$next  = \$signal$241 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          \$signal$241$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$241$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$242$next  = \$signal$242 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          \$signal$242$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$242$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$246$next  = \$signal$246 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          \$signal$246$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$246$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$247$next  = \$signal$247 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          \$signal$247$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$247$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$251$next  = \$signal$251 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          \$signal$251$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$251$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$252$next  = \$signal$252 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          \$signal$252$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$252$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$256$next  = \$signal$256 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          \$signal$256$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$256$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$257$next  = \$signal$257 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          \$signal$257$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$257$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$261$next  = \$signal$261 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          \$signal$261$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$261$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$85$next  = \$88 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$85$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$262$next  = \$signal$262 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          \$signal$262$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$262$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$266$next  = \$signal$266 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          \$signal$266$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$266$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$267$next  = \$signal$267 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          \$signal$267$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$267$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$271$next  = \$signal$271 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          \$signal$271$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$271$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$272$next  = \$signal$272 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          \$signal$272$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$272$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$276$next  = \$signal$276 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          \$signal$276$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$276$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$277$next  = \$signal$277 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          \$signal$277$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$277$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$281$next  = \$signal$281 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          \$signal$281$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$281$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$282$next  = \$signal$282 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          \$signal$282$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$282$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$286$next  = \$signal$286 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          \$signal$286$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$286$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$90$next  = \$93 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$90$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$287$next  = \$signal$287 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          \$signal$287$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$287$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$291$next  = \$signal$291 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd185:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd58:
          \$signal$291$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$291$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$292$next  = \$signal$292 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd185:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd58:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd122:
          \$signal$292$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$292$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$296$next  = \$signal$296 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd185:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd58:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd122:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd186:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd59:
          \$signal$296$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$296$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$297$next  = \$signal$297 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd185:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd58:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd122:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd186:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd59:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd123:
          \$signal$297$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$297$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$301$next  = \$signal$301 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd185:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd58:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd122:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd186:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd59:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd123:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd187:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd60:
          \$signal$301$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$301$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$302$next  = \$signal$302 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd185:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd58:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd122:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd186:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd59:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd123:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd187:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd60:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd124:
          \$signal$302$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$302$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$306$next  = \$signal$306 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd185:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd58:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd122:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd186:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd59:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd123:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd187:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd60:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd124:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd188:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd61:
          \$signal$306$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$306$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$307$next  = \$signal$307 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd185:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd58:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd122:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd186:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd59:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd123:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd187:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd60:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd124:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd188:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd61:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd125:
          \$signal$307$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$307$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$311$next  = \$signal$311 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd185:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd58:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd122:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd186:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd59:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd123:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd187:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd60:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd124:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd188:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd61:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd125:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd189:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd62:
          \$signal$311$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$311$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$95$next  = \$98 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$95$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$312$next  = \$signal$312 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd185:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd58:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd122:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd186:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd59:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd123:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd187:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd60:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd124:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd188:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd61:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd125:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd189:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd62:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd126:
          \$signal$312$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$312$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$316$next  = \$signal$316 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd185:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd58:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd122:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd186:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd59:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd123:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd187:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd60:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd124:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd188:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd61:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd125:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd189:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd62:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd126:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd190:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd63:
          \$signal$316$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$316$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$317$next  = \$signal$317 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd185:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd58:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd122:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd186:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd59:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd123:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd187:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd60:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd124:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd188:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd61:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd125:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd189:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd62:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd126:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd190:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd63:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd127:
          \$signal$317$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$317$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \ack$next  = ack;
    (* src = "/home/james/systolicArray.py:34" *)
    casez (\$320 )
      /* src = "/home/james/systolicArray.py:34" */
      1'h1:
          \ack$next  = 1'h1;
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \ack$next  = 1'h0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$10$next  = \$13 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$10$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$100$next  = \$103 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$100$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$105$next  = \$108 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$105$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$110$next  = \$113 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$110$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$115$next  = \$118 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$115$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$120$next  = \$123 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$120$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$125$next  = \$128 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$125$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$130$next  = \$133 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$130$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$135$next  = \$138 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$135$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$140$next  = \$143 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$140$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$145$next  = \$148 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$145$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$15$next  = \$18 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$15$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$150$next  = \$153 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$150$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$155$next  = \$158 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$155$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$160$next  = \$163 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$160$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$165$next  = \$168 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$165$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$170$next  = \$173 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$170$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$175$next  = \$178 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$175$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$180$next  = \$183 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$180$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$185$next  = \$188 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$185$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$190$next  = \$193 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$190$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$195$next  = \$198 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$195$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$20$next  = \$23 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$20$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$200$next  = \$203 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$200$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$205$next  = \$208 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$205$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$210$next  = \$213 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$210$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$215$next  = \$218 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$215$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$220$next  = \$223 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$220$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$225$next  = \$228 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$225$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$230$next  = \$233 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$230$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$235$next  = \$238 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$235$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$240$next  = \$243 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$240$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$245$next  = \$248 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$245$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$25$next  = \$28 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$25$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$250$next  = \$253 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$250$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$255$next  = \$258 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$255$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$260$next  = \$263 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$260$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$265$next  = \$268 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$265$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$270$next  = \$273 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$270$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$275$next  = \$278 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$275$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$280$next  = \$283 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$280$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$285$next  = \$288 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$285$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$290$next  = \$293 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$290$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$295$next  = \$298 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$295$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$30$next  = \$33 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$30$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$300$next  = \$303 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$300$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$305$next  = \$308 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$305$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$310$next  = \$313 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$310$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$315$next  = \$318 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$315$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$1$next  = \$signal$1 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          \$signal$1$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$1$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$2$next  = \$signal$2 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          \$signal$2$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$2$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    dat_r = 32'd0;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          dat_r = \$signal ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          dat_r = \$signal$5 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          dat_r = \$signal$10 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          dat_r = \$signal$15 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          dat_r = \$signal$20 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          dat_r = \$signal$25 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          dat_r = \$signal$30 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          dat_r = \$signal$35 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          dat_r = \$signal$40 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          dat_r = \$signal$45 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          dat_r = \$signal$50 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          dat_r = \$signal$55 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          dat_r = \$signal$60 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          dat_r = \$signal$65 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          dat_r = \$signal$70 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          dat_r = \$signal$75 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          dat_r = \$signal$80 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd81:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd145:
          dat_r = \$signal$85 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd18:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd82:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd146:
          dat_r = \$signal$90 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd19:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd83:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd147:
          dat_r = \$signal$95 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd20:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd84:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd148:
          dat_r = \$signal$100 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd21:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd85:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd149:
          dat_r = \$signal$105 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd22:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd86:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd150:
          dat_r = \$signal$110 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd23:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd87:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd151:
          dat_r = \$signal$115 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd24:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd88:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd152:
          dat_r = \$signal$120 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd25:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd89:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd153:
          dat_r = \$signal$125 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd26:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd90:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd154:
          dat_r = \$signal$130 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd27:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd91:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd155:
          dat_r = \$signal$135 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd28:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd92:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd156:
          dat_r = \$signal$140 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd29:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd93:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd157:
          dat_r = \$signal$145 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd30:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd94:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd158:
          dat_r = \$signal$150 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd31:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd95:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd159:
          dat_r = \$signal$155 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd32:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd96:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd160:
          dat_r = \$signal$160 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd33:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd97:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd161:
          dat_r = \$signal$165 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd34:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd98:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd162:
          dat_r = \$signal$170 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd35:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd99:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd163:
          dat_r = \$signal$175 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd36:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd100:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd164:
          dat_r = \$signal$180 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd37:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd101:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd165:
          dat_r = \$signal$185 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd38:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd102:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd166:
          dat_r = \$signal$190 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd39:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd103:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd167:
          dat_r = \$signal$195 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd40:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd104:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd168:
          dat_r = \$signal$200 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd41:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd105:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd169:
          dat_r = \$signal$205 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd42:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd106:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd170:
          dat_r = \$signal$210 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd43:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd107:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd171:
          dat_r = \$signal$215 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd44:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd108:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd172:
          dat_r = \$signal$220 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd45:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd109:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd173:
          dat_r = \$signal$225 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd46:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd110:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd174:
          dat_r = \$signal$230 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd47:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd111:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd175:
          dat_r = \$signal$235 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd48:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd112:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd176:
          dat_r = \$signal$240 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd49:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd113:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd177:
          dat_r = \$signal$245 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd50:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd114:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd178:
          dat_r = \$signal$250 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd51:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd115:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd179:
          dat_r = \$signal$255 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd52:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd116:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd180:
          dat_r = \$signal$260 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd53:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd117:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd181:
          dat_r = \$signal$265 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd54:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd118:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd182:
          dat_r = \$signal$270 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd55:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd119:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd183:
          dat_r = \$signal$275 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd56:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd120:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd184:
          dat_r = \$signal$280 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd57:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd121:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd185:
          dat_r = \$signal$285 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd58:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd122:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd186:
          dat_r = \$signal$290 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd59:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd123:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd187:
          dat_r = \$signal$295 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd60:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd124:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd188:
          dat_r = \$signal$300 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd61:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd125:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd189:
          dat_r = \$signal$305 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd62:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd126:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd190:
          dat_r = \$signal$310 ;
      /* src = "/home/james/systolicArray.py:26" */
      32'd63:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd127:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd191:
          dat_r = \$signal$315 ;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$6$next  = \$signal$6 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          \$signal$6$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$6$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$7$next  = \$signal$7 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          \$signal$7$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$7$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$11$next  = \$signal$11 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          \$signal$11$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$11$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$35$next  = \$38 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$35$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$12$next  = \$signal$12 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          \$signal$12$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$12$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$16$next  = \$signal$16 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          \$signal$16$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$16$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$17$next  = \$signal$17 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          \$signal$17$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$17$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$21$next  = \$signal$21 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          \$signal$21$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$21$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$22$next  = \$signal$22 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          \$signal$22$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$22$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$26$next  = \$signal$26 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          \$signal$26$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$26$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$27$next  = \$signal$27 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          \$signal$27$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$27$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$31$next  = \$signal$31 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          \$signal$31$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$31$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$32$next  = \$signal$32 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          \$signal$32$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$32$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$36$next  = \$signal$36 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          \$signal$36$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$36$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$40$next  = \$43 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$40$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$37$next  = \$signal$37 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          \$signal$37$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$37$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$41$next  = \$signal$41 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          \$signal$41$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$41$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$42$next  = \$signal$42 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          \$signal$42$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$42$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$46$next  = \$signal$46 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          \$signal$46$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$46$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$47$next  = \$signal$47 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          \$signal$47$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$47$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$51$next  = \$signal$51 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          \$signal$51$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$51$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$52$next  = \$signal$52 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          \$signal$52$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$52$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$56$next  = \$signal$56 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          \$signal$56$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$56$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$57$next  = \$signal$57 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          \$signal$57$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$57$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$61$next  = \$signal$61 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          \$signal$61$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$61$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$45$next  = \$48 ;
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$45$next  = 32'd0;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$62$next  = \$signal$62 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          \$signal$62$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$62$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$66$next  = \$signal$66 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          \$signal$66$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$66$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$67$next  = \$signal$67 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          \$signal$67$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$67$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$71$next  = \$signal$71 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          \$signal$71$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$71$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$72$next  = \$signal$72 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          \$signal$72$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$72$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$76$next  = \$signal$76 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          \$signal$76$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$76$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$77$next  = \$signal$77 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          \$signal$77$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$77$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$81$next  = \$signal$81 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          \$signal$81$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$81$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$82$next  = \$signal$82 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          \$signal$82$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$82$next  = 16'h0000;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2097:dump_module$1 ) begin end
    \$signal$86$next  = \$signal$86 ;
    (* src = "/home/james/systolicArray.py:24" *)
    casez (adr)
      /* src = "/home/james/systolicArray.py:26" */
      32'd0:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd64:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd128:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd1:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd65:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd129:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd2:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd66:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd130:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd3:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd67:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd131:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd4:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd68:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd132:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd5:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd69:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd133:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd6:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd70:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd134:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd7:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd71:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd135:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd8:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd72:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd136:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd9:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd73:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd137:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd10:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd74:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd138:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd11:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd75:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd139:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd12:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd76:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd140:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd13:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd77:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd141:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd14:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd78:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd142:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd15:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd79:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd143:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd16:
          /* empty */;
      /* src = "/home/james/systolicArray.py:28" */
      32'd80:
          /* empty */;
      /* src = "/home/james/systolicArray.py:30" */
      32'd144:
          /* empty */;
      /* src = "/home/james/systolicArray.py:26" */
      32'd17:
          \$signal$86$next  = dat_w[15:0];
    endcase
    (* src = "/home/james/.local/lib/python3.10/site-packages/amaranth/hdl/xfrm.py:503" *)
    casez (rst)
      1'h1:
          \$signal$86$next  = 16'h0000;
    endcase
  end
endmodule


`default_nettype wire